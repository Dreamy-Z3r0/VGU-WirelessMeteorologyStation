** Profile: "SCHEMATIC1-freq_response"  [ H:\OneDrive\Senior Project & Bachelor Thesis\Personal works\VGU-WirelessMeteorologyStation\01 - Simulations\Archive - from Senior Project\LPF\Analog RC Filter\01-ChebyshevLPF\chebyshevlpf-pspicefiles\schematic1\freq_response.sim ] 

** Creating circuit file "freq_response.cir" 
** WARNING: THIS AUTOMATICALLY GENERATED FILE MAY BE OVERWRITTEN BY SUBSEQUENT SIMULATIONS

*Libraries: 
* Profile Libraries :
* Local Libraries :
* From [PSPICE NETLIST] section of C:\Users\Z3r0\AppData\Roaming\SPB_Data\cdssetup\OrCAD_PSpice/16.6.0/PSpice.ini file:
.lib "nom.lib" 

*Analysis directives: 
.AC LIN 100 10 120Meg
.OPTIONS ADVCONV
.PROBE64 V(alias(*)) I(alias(*)) W(alias(*)) D(alias(*)) NOISE(alias(*)) 
.INC "..\SCHEMATIC1.net" 


.END
